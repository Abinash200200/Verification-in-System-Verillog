class trans;    // Class declaration
  bit t;        // Declare a bit type variable 't'
  reg q;        // Declare a reg type variable 'q'
  bit clk;      // Declare a bit type variable 'clk'
  bit reset;    // Declare a bit type variable 'reset'
endclass        // End of class declaration
