interface inter;
  
  logic clk;    // Clock signal
  logic reset;  // Reset signal
  logic t;      // T (toggle) input signal
  logic q;      // Output signal

endinterface
